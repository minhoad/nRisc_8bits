library verilog;
use verilog.vl_types.all;
entity registers_bank_simulation is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic
    );
end registers_bank_simulation;
