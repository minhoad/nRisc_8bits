library verilog;
use verilog.vl_types.all;
entity ula_simulation is
    port(
        a               : in     vl_logic;
        b               : out    vl_logic
    );
end ula_simulation;
