library verilog;
use verilog.vl_types.all;
entity pc_simulation is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic
    );
end pc_simulation;
