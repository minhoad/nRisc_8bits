library verilog;
use verilog.vl_types.all;
entity extensor_de_sinal_simulation is
    port(
        a               : in     vl_logic;
        b               : out    vl_logic
    );
end extensor_de_sinal_simulation;
