library verilog;
use verilog.vl_types.all;
entity data_memory_simulation is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic
    );
end data_memory_simulation;
