library verilog;
use verilog.vl_types.all;
entity mux_simulation is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic
    );
end mux_simulation;
