library verilog;
use verilog.vl_types.all;
entity unidade_de_controle_simulation is
    port(
        a               : in     vl_logic;
        b               : out    vl_logic
    );
end unidade_de_controle_simulation;
